`include "includeme.svh"

module bottom (
    input  newtype_t a_i,
    output newtype_t y_o
);

    assign y_o = a_i;

endmodule
